`include "mips.v"

module test;
endmodule